package mem_env_pack;
`include "mem_sequence.sv"
`include "mem_scoreboard.sv"
`include "mem_subscriber.sv"
`include "mem_agent_1_sequencer.sv"
`include "mem_agent_1_driver.sv"
`include "mem_agent_1_monitor.sv"
`include "mem_agent_1.sv"
endpackage: mem_env_pack

