class mem_scoreboard;

    mem_sequence trans_sc_br;

endclass